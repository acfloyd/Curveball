
module Frame_Score(
	input clk,
	input rst,
	input[15:0] your_score,
	input[15:0] their_score,
	input[15:0] game_state,
	input[15:0] pixel_x,
	input[15:0] pixel_y,
	output[2:0] color
    );
	
endmodule
