

module Graphics_ASIC(
    input clk,
	input rst,
	input[3:0] chipselect,
	input[15:0] databus,
    output[23:0] color,
    output[18:0] address
    );
	
endmodule