
module Ball(
	input clk,
	input rst,
	input[15:0] x_loc,
	input[15:0] y_loc,
	input[15:0] z_loc,
	input[15:0] pixel_x,
	input[15:0] pixel_y,
	output[2:0] color
    );
	
endmodule
